entity MAE_emission is
	port();
end entity MAE_emission;